‌‌‌‌‌‌.include spice_lib/sky130.lib
.include PFD.spice

XX1 Ref_Clk Up Down Clk2 GND VDD PFD


v1 VDD GND 1.8
v2 Ref_Clk 0 PULSE 0 1.8 0n 6p 6p 40ns 80ns
v3 Clk2 0 PULSE 0 1.8 10n 6p 6p 40ns 80ns

.control
tran 0.1ns 5us
plot v(Ref_Clk)+4 v(Clk2)+2 v(Up) v(Down)+2
.endc

.end
